`define OP_LF       4'b0001
`define OP_LS       4'b0010
`define OP_LI       4'b0011
`define OP_DC       4'b0100

`define MEM_DELAY   7
